module pseudo_DRAM#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=128) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface
      // axi write address channel
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [7:0]             awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------

      // axi write data channel
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,

      // axi write response channel
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master
      input wire                  bready_s_inf,
      // -----------------------------

      // axi read address channel
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [7:0]             arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------

      // axi read data channel
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);

/* vvvvv  You can only modify the 2 lines below vvvvv */

parameter DRAM_p_r = "../00_TESTBED/DRAM/dram_0.dat";
parameter DRAM_R_LAT = 50, DRAM_W_LAT = 50, MAX_WAIT_READY_CYCLE = 300;

/* ^^^^^  You can only modify the 2 lines above ^^^^^ */

//  --------------------------------------- READ ME ---------------------------------------
//
// Modify your "dat" in this directory path to initialized DRAM Value
// Modify DRAM_R_LAT           for Initial Read Data Latency,
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//  ----------------------------------------------------------------------------------------


reg	[7:0]	DRAM_r	[0:327679];   // addr from 00000000 to 0004FFFF
integer dram_r_lat = DRAM_R_LAT;
integer dram_w_lat = DRAM_W_LAT;
//--------------- encrypted from here ---------------

//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
cCr3WnORX7ZoR2xgRWHsUnlYx5MnfAyA9eiWkuoIlx76GFXPvlF+XAA2JBBCuKO/
wJeXSB7AtRSeNC8sSQnIS0Fc9yAbDmOaBhGRAS/1Vm2acsmX5v+YeHXB831qYi7s
Ra8yj0KmoafhJiycvhP3ZtBLRdDhZ45pgDrKjt4RxcF8fBVDLE+fc4rh+6s8NkK2
HSJZcPop+tAOMacQq0nh1TbtBux952Y9rBiSvp/zwJRxHEY2i2U9biVvnBAJ1nqu
HjuE/hNrm7hKmHpXCYT94t59+Zwvbz0+6ZB8m0DzA8V7PVpH4mrIQmzS79zsskV6
4eHU5ODj6uAJ+mDG2dv36A==
//pragma protect end_key_block
//pragma protect digest_block
o/0i2xv1q0UkfQbWtgbvEMUzraM=
//pragma protect end_digest_block
//pragma protect data_block
2kixBNchFCR+YxgV6251+qONuf96NvnrH0a4fqv0dMQf80HwinlkxgmS+JcLrpYS
GyvD/6BdJADJh4XApftIG09Y7M9nB+9yUxq9y3H5f3FiclkNezpRCYOpdKgIPpD2
+DcoNTW1cqbrEi449zo0ZRvTHDsi7RJdZJJQ/5vx7khjKdXIYjvWu1/BGS8BduJQ
bE2tkAf4UoiIYjm+d3Ot7owK8LcEetG/RVO0fwT9GQavVBB7PSA+zynqtMUM08bk
BTRgrQAJnyK0xpVllwNALv7IfBL3xBKHSflQyGhmW4t5EzqJby8jXFQOpcoNV4M7
o+lo0Ak8Yeg5e+DKlXi9aBPy0EwJHebTgk3Z0dC/A9FULx2cLjc+R499rqispUmC
6fpUp4WNwrZgXYObSadAZYvup7UrEU1bMwswKReO/Ep+wMv/hlZFyEExxFK2l5wN
IS3imCnyW94U9+qJs3r6xeJr+Dl+tLnyF7rKk8QSso70OAQdvprPzI/QsTfr6C0e
I3BTJnnE1EnUrps87/64UcJB/YzTMUudol3UejEA6Lge/OsVF57/nHohSybWnZJg
zEcCxt7ddzrjtb1JarbYenRhODqar3pYI4KhaVVu9OsQ0bfPyFj0FaUZ40dgiRKI
bPDAU1unMxWKsrVr/cNA7b9t1MBWen2/h/9UEf0ztJEmeMhQ6v3QkVTTfh+YHoSm
6k8PFuCVm6dH1AppQ6WObs78eHr9OwqRGq49Mbt+h11FRYhNh0t2gvRHzYS4670d
G7QlffC/cDI9tPx3d0vIok6196XrdZr9Ta349HlK7Kwtg0kPYmN8/27SuolmliTI
4cZ1DJFYB7sErCAfXYXiMvMEMUt72QWqy9fao2wMb6f/+/4rS/1AYUTu0fkOqCuj
saXccA6s4aKZ9aeo1x6Hx472hXVr2agYtNSjG3UzGnk2oOxNjnkVLUfHRJsBBD7j
08ioEvOYBWw5NK7lx6uWyCt4/polVSz2e1UzvVsPzz0DO8Dyb3C88hUz0G3sUDTz
hgSthcUZtGzWtEjCOA5d1VvLq86Rl5d3xC3QrN83foijfpLebyeNzx4qqEaN6tie
t0uVuS6o8j0mmjaJIfJ+vu0Cvp7eJ18lozmhfh3A9C7JfwC9oy6OpGq22HdbcXo7
tDyePdJy3DtEpVoPQ9/RxCBaJVsFa04aPRCUpguBtfhCAoPpkomtqlJOsq+2uf6O
juGU8CfuW8zQVskjf3VBLkgeLZ55M3wcpDJFtp0laYB3V/LxrO5ik+qhK2I/f+80
yXDSv/nTeFEjUhzMysfZj0FF9BUaNvJBkj94lqW2Da7opTa6N0Kn4M6HJY2DDzYY
VoKwtvLrQzd6awZsXyBTPc2ZKE8AD7opR3uFD1cn+m82vk+QtIP4FkC40Ne4Gsrj
fkxcLGxA6lUJOrDgxnIcjyaKQ1QErr9Mdi91UFEJ+6QnFL6Yl2vu67507cECxtI6
KtRlHk0TrEeOr5T+2el/LxlKjmudn0uyeW0Hm2eA8U/kxwDNv8YJcpmTWjOGQY64
sJ2AnQQQra9hqxbugj+fZ1fdZgKRvIKhBjAcZ8Gl6PFxkrcDmJEHv9mvJiVRT9Wl
4wCkIWi6b2A/fcDGuzzcasrevmuhOM/LjjomgC5RUms6sY2JgNzz13a4JhmpSKgG
hc/QsYCGmq9zKVi+8Ws9+QM0b8LEUN4RzG3jN2/0JgwEj//a89lXJZNhL6fLtQOa
yxKKr+XNTKKJ4ewIK1xbj5+PP+QcYZ6Qm4d/FLuFvzC6970yhFoXFN9aT9tTjGzP
V9qzc8VbTIQZDLsp7j2inx/vD8vTOc/75K0lhaOTXIIBQJ++M8HX/DltYhu2S8Qx
itg6J9iv04rub0ASPYJ5tbOgjotBwd6AZChVz5WPLNsEsMk2Ge7BXex8T756JoQ9
2o5lF7ePW9PEp3sJd3W4xF/Dnfv5tUy4jLQwJZ+5BBQcqm4oNb+nTake/7cPxoYj
C4Qq6se9V+GNsslzqb7k2XqqEGWtMH6Ypb5CQqzFtQtmDX+zwetReZw++0MChWPM
iqbLjdqJPg6d2YC4GPcnIsIuxulaWFrF3kKEFHVFsO7t7ZfSQXtbJV0j6Ztkxtf4
pnkt19g+Bn46L8Jbl5C32b8tXeiKQSRtqTdN9LQ7vAhtzGcI8jhQj/38jGJZgWKy
bPIyC71P3S79D8fTbbLfH5MoVs468nk+Jlpy7s9mNzwJrsO2MhehQlqXOpM9GemZ
cBPjDFIvr+TwqY+WifiadaZyJU+s9fuToG1Mi/QKMxwggUTZXyN7qd8OsIfKKWfL
2W7kesU0LZBHqko9N5sjA06Bj/nqUnZgjFFRMn9KU7Zh7ZO3SFpz6TIO3OYID8cJ
MO3sPZ/fq2Is6k/SQ0R11DWeKxn1auJv3A90LP3wmUalGO7ofQvnhX+9ScT+eyAJ
1SmWqMw8G+w1osMqIdnlE+E+iFcgWuw6DZfIqwU/tTwcYs95L9HHMk66lH+oW2fr
ywEub2wG631f5XJsMl4XaRFvO3XjFENbR4IiDZ72QbL9jFRQf7sekANV2lQ1u6hT
JLNCOrv7CN4bDlZWYU2z16ua5PCaJYvYaeYFWpyfOAEUJJJaj6mBc4KQuAAmZ7H4
vD3ENre224idkz47SJ5BarnaR39csCyaZxuW/v8Nk7uReTSdru7LBiLfHoGg0PbN
AskS2UAmg7Ps9ET3jBYlv9pcfxJR4bXXgK5rYeZHiHT57SlBtHzb5oNVklVZi2AG
PO+x+gF4MAPlj62fscai3UprrBSKEkfMfSgO77MIxKAW9h3ik4RlFJ6jnDIHtf9l
l2xIAidcE8uBy+WuC0TjNE75kBWI2n51RMzvW7WUeRcuiUae0LOtzcD0Aqx6k8Te
t8dJYEKgpf8/0O3OU3fKPwvXg6RgSOuQZgtiEyDeJzDfCZqd6vz7ewVGxmPxtXwC
O36dfqcb5QgmMbRwYFLDmgSzgxn6yCRe+odGQi2tGJ4wpQbcoWyIUP5ZF4ZPfk0l
uzKxakkOoL5d5UhlEyizhfRRAM+IxuEfzfByP2BE6zLkanTNDiVrG1RoV3/a/YLh
dVcjOu+gdOaALd/7lCBxpvyXsYtvISX5Vem/VgM3VXM1raVWBeVkjApXuxBqJvpa
oF3e8gMCZr/wVK8eS+WziUAHvuRRNsEufNd/VTQQCL7QZKMz9h8dza7ZEvep9o/m
mktwyv+LP4LK3A3xpgcW/AUoayjr/agd7HvL47/1WOh0Czt+KOMCERrgwb+4mZ+K
SJRtyaqSqZ9iAZEMiaNiBHa5Qa5pOqZEeoZ5A/zQ6xvjLFmEzlI7vOyH6iRoeoiq
RDXe/molnk8JYF3ZDsCOoWZY5MKOKqLtxv67AUBpMmNgkozGqvFnENa2uKxmFVNO
PjUt0GFb4C0qT35e3OcWi0PvRy3A3UsTxoVCJAyoe2UNHAMlSXMZ85pjsuJ5tQmI
P6UfiEjHZ6NC5QijEDFz4mL9N9F8ATyhHt0NCX73Ibykrei+Vn0UgzBb9BXhkACZ
Gy1ONBXx22CDgv4pUer+eEJS1AcasHth46U7AVmFEAwaXztDQGclGOBgFOzuAmzi
p/D9NsYehnDLO3KMIVJAPQOeftukA6Eb0u7iA5r1QQvRs/9OSiLvY14XbRukvGQm
TLdfVDVV6FQyxoKll3yJw6FVP6v1gsH/9uCZ7EYKoK3dxrKRMy+qdbdhQ7Ccch7K
pij7rggCPJsthwWPLHCcLDiSsifvV205R/yeBdppxKksGEJDzWNquAwr630WOVpI
12o02ORt4/mqppswXofTqfbN8mKg468l6IMArxVhDii9FpKf6ICXW8/e0Arz0mxB
xxoGkzyFeOF6ECKCL8D+lxZKIxA4VkcxDdYGGKuKYKZAiFDmRZ76QT/LBVUhM6hB
Y87a0kqdV7skZ4ddcCK9M0Qx3Tn53S4D0L6weSRTUEr4YhiHwyElaO+HNthaBH8O
rM3mcpRNiEpMwDpiq74lhw2YdnwdAjalwOmSeBrVxS+WRiJm90OnCsqwkYo2GyR0
+zJCJHgG/SPqqlLT0MU3kTAkmMMddVrJtAK6QQClG1Gw1RNrad67j3HdzeCjxSqT
yvKOlPSiMuzX6dyiLoK5CkhgBnlg9XjYjI9F4FLNdNm+29+iaPa76LDeasOrJmY+
E4xY+k+s1lCiQN/i8xLtv2MNN+y0amARdSjGB/JKZB7w9oIhc3QGu8idisVzjr5b
8UvlspSs4SIypwpcQCqIUGS2pMsM2nWIGbdsPGw9f9tj0IDm16Qs9wGSgEftWZ7P
6WPYNoXxy7cL8lJmww9AYbhF3C8Wp+1NQzAl1vsBpQqStCmXjluc+Qo4sdjRYX9m
le4RLLYo3nAO6AYqkCo0EGdLnxLAdgSMwoo90gHp3b5kqIp06AKWLBZz+NaOJJGT
FnqEECCqEO55XyF6mky36c9ON3v0LiMXdy1SGd9YmKiIxaIPwT1h0kIaTFWWTbMe
/nAl03fnElwMuE62ExhdyzmWEdSRhqI4WElbaanqKQ9WqZucXtoGjpqHwJpB6IuQ
HPjt2rfqAeG6LnuLkL2LNtrJ0OaoEFbtA4u+kRyVMeTZea/LabgARZX+wrfn6dZa
FqkiIn3PzIK5+JtvWnvaZEYmaAlmd26PIxcEivSJP0pGR/YIt1yFBo/X7rT7jbvn
ePIn91nJhGaETt3+LsVhFGk4E9ODUYIo7DgicdA5H/EgqepsXweEjlSTn70EOoZj
sbTVQiB05lK3jmtm6pLsDsl4NQzgi88wz4bgRu4K+2YQtIkTgo9gpFAHvl79vyhb
rvwVf/dJ+owjpmn0LrCti3EnJkBNO6pPlqh9T8qnEER1AXqpQ94+jQqAqSFbcrVm
Q6XGZkouH73OSMJZQApfAdQX9AB6uQ5rgfrWm2eu+qNHcDJHQ/LjaMxTVgFMkEP1
swLczttqRlcjJl1sH3LtaNX1zBA/qYSWXpItvPGPWCXmQiD3F6nk5zNy2tOChIaX
aVUhsgW/8ifnzYXMbhgYNe7bwcY34yoHkT1G6x49WEGDtqO53rz1m7zN5lEm2+op
JNqCiO34Ri42Be9OeDpO/AZg6xVTf2Gez7l3IphE0P1mqzcH9piWrDZocUcP7oYr
/4vEAzmdDN5I6wQz5YieBDS1dhCaqfvZF/P16HvgkoA3Mw13tgjTnm1QVnGBNY3p
c8Vhhsb1NyUF4Fpkmc4hwWg6j8r9X4syTVfT9zSfgj0Fx3HFUYzVvcqZTuhwiI9a
j7WpbxZBUkmYLuRRct3vHs3wUswBWY53Phpbn5e3D7MWlpAXhsfa9/9JqEcH1wrR
4JdSHNkulpYbIZp3owRzcJ/s+8mkjc+egWL+M4UFGxGgoPQKZretDYBrdiehBVR4
Nmm8szOWYSOBQWoxPGzUuSqSkUaE13jj7yG4/nvuNcIS6H0bawj0KdGfRGSnsVHL
eXMoTI1//evDVkgESS5VvsD01J/bqYz+ZzjPcS4QqYW/BI+uOSnG6Jpd45kxPw8h
m1nbqLNw4NXonfeuejDoY1TuqIyIOuGDDmBJNKGsxlEZvCClqL1bGbMMYv0RJM3G
FRzToyNvn14rA1w7GdgUtdlN4fC8/5leqXBWRBtiyODNB6wtAnaR1nG5IK95XGiU
YnrqQaeVsuldTZQ5MBAekLpoRr+VnlzpX9d2EBxLrdeVc/X/wHcyEu/RDOSMk9Wu
1+3+udMv8uP+xqrBzykG6fBkZG2womySWzU1oXXxYHgIQoX6b4WBpUcEpBjfbb2f
sxUo/tnU4t2DrXhSir1xVXbPDVUY0LxnHZrRAvldxIOOKvB+IXkqRPO+bzwVVHBa
WnTIsLTbMwnucBh4J5inGPi0RXPYSEw6l2RsQmaWMxa4zyKvYGiI4tIc/Sat56WR
zuAIiKa9eYW9LcR8qCeFRcguzM6F/2CB/+80FatG1rEVemNfc/vnzwskyuzmD0U0
3FJN1hinqE4q/iN8WOmuO/dFiuDGZrSgAYRvV/wI8fA89jKErVOnXVJxPd6Colcp
E6LRlIZ+E8wxcr9rKzX9n1uT85h8JN0wcwUKv/e2qa2kDdq5Y07/bObLu49KVYrF
n3iGB/uOtJyQUU3TEY1WM1wOqiY8/DIEcBpUkDkZZgy1e78qUVzhWqFKDQUqvwHI
5bTuUf+GeRl+dYsyZI4CUg8tm6KhjYs2qoKkUBQ2HiwJaftdboADjF2+92vtQnu6
7/g6G9DyeyASpZHfohgDdQZIeQprtQYcvq5+DpG64IzNs3oaZucU54GSahBqn1pZ
ll6fLsN/XSGRRMZ5wkwoY6zRXHaSEsUr/ayqlzV0tA+oIfZZZpc/7zEubFq1A2Jg
nnEZT/44v3e2kXJDld9idZ0ZV7iO63noyr33sd+MkcYKDO34HJVtOkU8mrYjSp67
Dn050fbiQpA6+8bjmed1BEYaq1faADYya5rTWVYaifSRT4hK3LXKuwIfUep/PSyr
avn4Wje2gqSG842VPtht+a44ekkB/RB/WazJYn39wdzO/Zg2ERhvG27NbBwKYkkt
fVK3ZsBzE/RrlhWOLyviX5uQDspyp+UxBen6LR2Sy4l1DzRYSK6GfGcut6mi4hpc
0wc08lGKQVP+2MqoGvVj13IolMIsc92THQU9wGZQvTON+ML0f2WdpcYr5KsuqEaS
CLW98EY2gr1eT/4HZcvzDBawrn8p5lHjgdbpx1ATEU0jvuCRJIlhMekrKPteYLvP
Qq3Ln4rAeEfJwe1qyHgKSS6mX9MLx4MxrustrU4yDepEoKJxvhK92nCrki34sS2z
pKIJgwXVgftCnKX90sENjNP/Se7QRsZNAWs7RRX8lVBXa06qg+P3qcqX8V4POpch
dY2hYA8GtZ/J+up6x1UiHtllZffYbj2QhAleFxdgfSkFy1qXLPaLTa3Fhy+WCLpo
bhsNUh2jW94l/r/3sq+UCP6//Py38dTCVj37K4LDigw4IYiLw0N5cjBYPmTBupI7
iVC0Ei1EJMVzKoF7WJXKYD6iRMc3gcg0zZ0h51fJRP8+Yyp8bq4OwdW5+CFh9uMQ
RBT96KobpVYeRRVkom2FYgvaczw3o6pZR9PHSSpCPSVXc4brOiI2+8AVTb091xRU
W2tC6YG1N4Fl1sBF0O23HhimNi8nFBR4PMHT/FfaAHC2bhrSE5i79fIL/9jfEmin
HGtk3/pamU1T1RjSiUoelX7O5D0kp2d6xntwKsaOYHLKruEe/k/JY0Ayqc11Mmm0
Q6XlU/RJrQ9mFKmZHCe85w3MX1wC4bD9LA7PNJzm+sETZeWc4krSNsWl3WU+hDVU
idGD30gYfEi6sm3VELOx1v1sctDnC3se7z+rAlMLn1lUXIuEQQSPfUjRwcKQvaAU
/gbvzWXsNbCYXy4QTOOHhM8SJD+P8oc3Bd0hCV31k7D0VrykTT5tNMPxUQSXoKhd
7lmXcyYVO1hJqh3F16XvC5aUTb26RpVu30JuOm1JWgyaHihGZuWDFq8ZgOmhinIe
ye4j/kpaIGc5w2t522QliR/o3wUNMIQNWOocSbj7ltAASSXHw63SfsA2dMjZonQQ
k5XrDbKRfAL13XQMAfw6qy/vzvaagNyxKKkwUE3Fubb0JO+AoY7uwsz33U52dNkk
sKVNybMf/s6xF4jbLyu/O4Re8p/8le7Ei4lqEr3EMysqfShNHzZuwtCVFbAPzqPh
kA5a8pyolml9GwzcZcCGCgmyKxzt47pAzUskUfjoTeYwufScXuBwwMYXhcIwUBLA
lhJq9PBo7CYxuCjG8Bs7hh6hL4kHZtOGcw82r651qNmJ+VNap8C3eM1tJShY7HB4
ftUUUNPVcFL+0Nmd4lRi/qUbyFwAOJ1OSbYxLGpKE58Au0KcOWRSsyZK9ye8O25O
IWK0ySHOWmo2KzWdkwh3pjuLWFMM8RYE7g4AzBVgpz7SnESWj4H4i5PnxmtERocx
fx4zk1wTAYv3h0LX0bC6rVySXj3XEa9lfdlv66j3X9adhpE5CrMuNQuzhUC8wJdh
gw7ELyOZdf2ybp56Bk+2ZMdvooXNoDUQNjgU6+V7zOlXna19FDLTOikybrQ0YFNd
HINBPJwR7QpS5sAc4e8xZ1NmCMQLIG3bH0hIY242KYjpJR3xdSvWp81XCGzS1o0C
1NQCatmshygsSGvzTjJyWc5TqPbbDML/boBP+9QCOl7S8OKsHocsyjY+OAK9Jc/N
jdE2jyeRtIhaLWe6uBNKcNcbitmBErjU/gIH2rDoG4yH9RCDaNMx46y2RbQ4OT2c
l4ATQB/kh0jPlqYJK8jW391+EZAEyZs7fE6RjShiggRKjQj0oXNC029IadQAZk/6
HNnx/TWRHCoOWy6jKcvbt3dZRI+R19QXJk7+n4Lsg/MstXiZeHO8QQgz0GozdbxZ
GnOeL+QSagMcSw1r5RXBOleahS0XXOFwEoff5AHovyA24zfVKVHm4U1gSFRGjQb5
Oy0DptIA6zNSBllSetxPTpFrEaPtw+9RpUO2BjLbijUW9V72adqWQPhZEpU6T0+h
ow1yV55d+x2Ih2DsTjVbCtX4mUo1li2G/Estqd5aGclxCFRznBdHqUY6J6OBkUpL
IYgdLDbgxkJFCyMqRqX8Hs7+aN/bkq+6EuRuU99vEkfhlwj7CsUtwfDCct7qf7VT
yquEtJNngFy2bMh9vIEpxcOOIJcTNw6dRnJsocwBcjoTcjEQ5bfB+iPIryLLRjIC
vJLNkhtseqBDArajCGT88Vs2Sqf35YAUDenqX+EOC1cjI8Y+q/p8uxK4aUoQfS1e
LjCXBcXtFQdSV3foqDzANs1W/gtmR6z0y5+pbTSULm0ADnya9XU8tBkc5EHhx9zy
r+MvFAtfhnEr1HewL+1xnQof8Gmth0RS51WaIFy7pEzRFo/d67ez36SGwWQgVdon
zKHgRCqKRNjEUCSQ3R5OzCPF5lJm14flh+/g7RGbZDArCxPxJjZwzyaJLdKPBqcV
XxSqG5KiMx8fDnFMUhk0ZEnEvGSJgprMhFPRDxCWaZMkO8+jNZHrHpDzGlPb7sS1
xMIljtoN/81Rg8cjpQqu/gO0U8s6NtOcMyIGinuLQHY4780NDkpn59FT/s/MVv22
uy0aaNBdU+GnTFI7U6TRKE6wJ6r6cxsvgqacbLDfM5LoB2lYPZT6QOBLlSK6yrj0
7aRBIQVlhGw6Rcs1Nh97dLVqL+NSOzV3o27QfmATmgWlg6wGRZXZibK45JU/nF8u
wNymqgEFjk/UjUnSirNMKlKt7+s9fx+d7lsS3gCakKTp7qqZ6k6Qd4ZyejFFys7n
IhTgWPnnPxz5J74UJ4hwbUyjJehXCJrmbyAnepGGjl2052ljfJ+SB5LrOaxnTc7W
x4078byW5ahPZ/CX2mc4C4y0CqApAEIM6w0UpD0ouZ+3M9VhTi6rDdDZoZ4aEaXk
IC4HBlOU7C0li6jZculPV+ZRcqKsaURZoVa+wqhCnEmQWvV1SES3VK72EGqcSyYa
oJHLSGDO7OP625McCSZdpBU9f4DrH7kr3Vn9s5/tuoiGu0Nd1dXCOWxJYEY4tEai
0MASfM9hziNG3HNBUWQGq+i8FC0oE/yKsxi0Tf6A4brDZKDl8+EQmzx5RXacje4Y
ovrbfkCh6njZkfepcIbac3BjHXoWSuov7w3/sdNL9KlH4EfpOuZ/1I9YnmXWnn9N
Eem89gDQqMisobj50ytEubSailotk/XzQCDJdSIZVtqkWauxG3YQFyqh/zilfBfV
Y4QO3e2g861XmpBWxzf4TqpYfx6/KjLCOfBrDKYtT8wswKZCpO8UpbnrGOGNcUdZ
DZTxw0AsMPN7VxLoMMgRwGtFi1Ez/6orblSgc3DhNWrzSvvNkKELnRfi0Idvi1GT
l1g7zHsmkjgQ6DhIP+wBIVDa1sMWCMesvLC49IPlhVnzHbN4dEJ+Po8nwrSAyrJF
8sq3vu7PD46teRqrVwzrgGMr/d64PjliDE9W2+1FbTl1TG8fHctbRgftjC9Saq9i
SsWO2AItlBwJ2kYpv9twI0Vxro8HrgLMSSom6PwZoWkEiQhuI9aMvX68lVuWtclk
t2xO6LSKfiGkXK+sPMdHiT0OMrcrxj2oTr0OEpGzgDvab8zGXMhl+rkatSdbcIGS
RF1Aj5Itsx/VdYKmDl9OA6p5ZJITBiLNCuXRj67p77b91kni+ytqBFqHPQDG8KDV
HeiasKYlyGKasc5Ps1qfDiTmh0VPVjaVcDgn5NI5Ypes8z9wAvZC+nPZtsuPYcrs
b1OBMnRurbCEO7z3INERsMQIHyv6A7LiHPBgY+ellE68S4cxSzX373JjyBeHhIHP
If+vcrBGQ9DE1IrzuWvFotiR2RluzN9N+CUweBctxWW8e75ny399CbWYspivVh6O
pcmpt846JkahnwRqAENcTjzbsxA4l95pOxJfn4cZ+6uc5xO1u8jrhrHa+KjvCMdL
dxf6k1ovTrH23AInlsqGWkUhVIZ3jGbYP/AwmgAAJcqdOXJvWQWLIhCSzJMYy+Tx
yNP2xgwEwOUpBS1PuS7z0mp24dXwYlG+qS+XQT/BStmlvlCoqjNQiBivkdBhTncK
Dkp4Fj6LIi6nAXsa1XXEQ5oR6/zf9CHTovOV2Klf6a84SXqlk3o6R456ociWjXC2
Z0p7BowNxBJ6w3H7QREGDxyQkZ5+gvPyGDeHGxtP6Yhz/oY9A9HxhfaTRB4tFEwv
wmJXwB4xHgBqQkfKNg0YPWq02w63nXSq3R4FnPRH5xNCCOwErNUniYWjQONRFSxq
scs5erCHSIzVnLpLmR0sWmMn1cHlGfsgq8JcIxb22PRH/9Ova6tslbeIktIbSuFE
HgyTQGEinl0Kl0O3kJwPzAxkL0VlnaCREJvijKHaHSS09lUV1QytdpvLr6S9RDnV
7BB/q6/6g00P/ynrdjr7P5U9O9T0R3ztpujsRH2D/L8EOdpliUsj2mAw2f0QtWa8
kCBC+wANuVbN+Rdhqka22JRa1vSkNxERjBgt6PCVrDQAGLLwbwMsyxSc0qIU2ecC
TsyYY/whhySsSwr8jS8UWwU9/lX56h4YRc6JDSrj4J3XGcGkw+71aOOE8AdSLorC
gG2xfII9w35wqH5xXoagAUpv9DjeQ1484wV7zK/kQqYPltqrRbhEwelshw9xupQP
V1A7Koz3EM93FCn1C8Kp8zqKYkaTBo+hJFmn8Cl/KM82TJA/7oVI59ACLxrSK5oz
FZjNHlXynvCuJytIK6qnz+uqvmrP2QRl1JPGG3DQrBDsZsqNde2y51l6VrcIKhI8
T7FqGfNuiY2uM6/Kmw9+3duQJXkpmWjSh6/cjwYGkATPhXwTwuZ47OYlcMpGHiIF
WWR8bm9NQWWpLWkVEDzwaR1EbztppTFyEDwbJ8V/ssiYsyicXuGWDmm593YLdqIY
V1qGbV+60rLq5K0E8d/saCLmzyW4RoPWOwJLBzTy8qsLkojaDIi26BKAkQknruEk
u3rIojyBhrKQW0AfTP88BcS9srAG4cy3A3dr3tPCgfZEmMRDykugE8txWOLemQZq
xefIzvO0a1+5U+0wSAEnpqFygKXOXTEBUn/lP6km6gCBRmYjMbtg586IkmYCVnL8
/s0MHz5a0MrXtJI3o7eDCr2DOfhbQ8dWeG06MEetkESdi4tl8OzcfONrFOGRCjdo
cwEQ/exEDnpzQKOPghINWztWb4NbaG6BDruuRmkkLHVN7kX8VVN/pYUrC+EUMDp2
z7tTtKFSg2rQXKRHOTVD9eeHy7KEmzXC3jfU86SLWrFiEiajwIX8AVUHmOpSjQ+S
nEHBsnAQWW9iyIOIAWtuCTQCa6upnFknEZ13RSHxVQmRMEh5uYj+HTqBRd8SN3Up
NaPAvs3pYTpH1w/b9EkNczHDbtpSuKIUqSbMqKnQ84QtdTF6Hqb6RRkH9bBmlhe9
TKFXlrZCGjgK5Fzy1wvS6hNgN334w9xSIf8rcYB+EYTk4EdkdBOJ32zNX7/oTu/W
XWzc5MddBn3whX8Zs9RPsxYllTfWVU5jTx5hgZgAG2VEjlHM8HLG90TGGD7fRZ9o
tsomf3Ph3tAe+keOk5AKG81Qy+irSXxyVkFq2fcyNQaC4BrTz1e8oSwPcqKl3L7i
eBl0bEvfRHieVFc913HZUmdZT4CAtRseWunBS8wHXPGWv2N8vtI5lZjf2Kmoz18w
UqwHp1v5wYNddyJ8ycQAoa0HMu4Onz/L4/FMsPBggoRawLc25WSOjAaIfdh4IGkK
MljZ1eiTTCSmbjTXVoBg5YT87xa/0xX+Rh1ifiz11RDgHqWzMPB5U+CuvTHSL8r+
fbIKQK0IHGg8Ado3Ll/aSAMem/45PEvp8YZHLP/7mOyXZlZmK7r85cNEt3aK23O3
h5J7MzlVOamgKvWSMUyFOzW90MefNfk+wnMNlq2kLmcCje5WnnJacdz3d36rj4uo
IOhM1611Lp/0KZJTXWmvB8jA9bTsifOSPLeAJLTAboeA46psSYXgp2jX0vYJfJ0X
eOblqvGcFpX+z4XLLtjtB4UzrXFiO710gA+w++t/Sxk1G83hxuZ7yri8DzjJHr8f
EUi7q3qb0WA71VPZdt1UWhqlnhlIVWUufHpl8dzu0Nvq9WJ2kyOQF1l4X0lt+JIL
BleSd023Ta8WqST99j0veWWgoHZliNOxVvrstXwao19hi28lFb+Zm1qseOf94HSr
/R/QOWf8C/JXn1cYLZ6t6gnVrBS7Q2lu/cYxdIzUmA7WvJO8orssdQ+QfUKikIAS
bMuq2ZyFuDvQAiRIDvGwgJr91VSYlvewDeA5SySqEtJ4TiFHh4MizXERM+guMbtb
AxxCV654WfVMivQcgbM7Ya6LcdXmoTZnpL4mYtyZcEAo32tNlB2HnGVbDuzHra0s
1NQtE8AZFFEjNhjAwrFdsfgK25Bz94JZQygwyunDemtyAGtNcdPS7BhmtsdvA7RW
bGJF86F2FhdJ9Y92h52ifEal+UDmUJGQ47O2OHKOk+kRVCcTD5Ysd8Lrnr8O6TzR
fBoYeGY5f2uAXEkMBhoCb/hHFuY93Vp603gUWD/t1WbL8/ldqWiD+PC8W8RYOZjv
OHbFu1yRyTrMg0GxPZK4uVZyw3cxpe7yvhdNsZyb4aAKCBREmmipK4oBQkSpScq/
U6C8jTeU3pHJ5tAMG8/GXVni0btCoFfOL9hTF261Vk6AQ72A12udd4L0tlaQ2N6O
M67nm/6w8wJi/hf7GbAuyQESltc2ewGbCDrSjuGJaNj5Q7hZU+/TNp9EzaAMdKvy
fKrDmMuhyBgTsJ60g1viFCQjNlwaoTVaQOpEQrGZyM5x++K+1lvIhyKYi52F+O/p
PDJ6C1HxTQycyAa1aVs4ZEvoec8YS2UfbTnzxOihw3tKrX4+DzSXlCxx+dbgL+KS
MlJLpoUkE+cfNJjkZ/1vFUMzOQOwcnzLQVbOJidbqLqhtkYqmWuYS46QF08Kwfbv
INJfZB/4m05l6bXyV/aVFNDymfOjVPPZKFiiBNWsY9aKOrpbX8DsvSGQQvZfXg4l
EizdmNBO04Vd/qQtP1i0AyK1tgcst9+b94eBHTTIt+sLun5aOmh2qT3w5AeQ2c/M
poY/Ll5+5LguPYREN8N+iJvOLRypzT4xkjFF34btbeh50GhvnLEnM6JqYQZDNi1o
Lp4tYeNIqSgf7WrD7WQxKsZwnSRbzrnxzumVvMX1MLY/fbpV4z3zsPe0+sxu249k
W8AePlIDOOm0QNZgAgWY5Z5pnh2NE2L05NC98G90dNj2a9Ya206FlpzFpiHEo/kl
m12tJhoswsK3FNI2nQYYa4y/yJ2/DR3elBCyGRlcW+pCy0H0/EXpaXELbj9SwGkP
z0I60DuKf3GNnySO0gSn85E6W3vHJhSqLiVk6ePVGMbFvyfOw69NH2LyHYkF/8/L
Sbdr0J/qq42sEifW/vaE0LgIWxRF80yy3/Q9BhTGHMAEedOZwcu26cynmTGkkkk2
Y55IxDszs/0aCywGMNgXTGH0nLikjxnon3BOGzTK2hjMWil4t3qWpiNT7svBYMA0
mlKm2IxJciQcoys+rxxFwqstMNS7ikgmutXub5tzJzTU8dLXInfcGIBzfmqegBXG
PfFCaN2BnPDRvuwhNvo1R2cdzJOt4W4nk8UTsJALnJUMz+eWXGg+iSqNeKS/+Myf
/sJOW9whijNbxR+boDBrSuk/ilxFDbGHvSa+zVLcnUyVuXhbHOyzK8y0csQP268I
pCVm6StIK1F2CKrPAprKWEpCwpRzwOm0wdzPQikWhrSLfvM692Kx6s/YJj4CSuKc
78Ank7N4k04qgKdbmZ0QmGl8rrsgrrw1SHgZ36GgYJaAH67nozWWofvK+qZGFiyr
fJ2iHgNlGrOy4PSg5OZGH9turjMNxzTzQrGmvQC1fkmMhK5rkDE3mjvOdUJUrnJ1
yoBqPBAmPuYgSvSl06/9a9RNmjIL9AVJqr4B/y/PZGSXMQb8eRmPHXVCq3/S9hhf
7T6unxf+0E9Z8AyOAzXJQcmL9XK34bQiusqRadIB6OASi00ycZvN9Ilg4HgJ0tsP
Um88n4k/wUJVh3Yr33AjNsl+gEVV95u0e6/sX/IO+78WsQed5QVckal/GNp/TUKx
W14Lc120jymk96eqf1njYCbZqyoC8rasN4hljQSSIUJ2VNIZS1eM7ueL+hVoW+uO
KuwFL3UPKqJSRpY7OJIYV4wsYLQH+5VCjDb/GtQfg/IHMEmSBDTwkS0Xe0bufvG5
P6S74w3wDe3hjtEKKnC4LzGM/8vNG5augr+pNfJtLbAeBw3/nprbj7NqZu8s2oOi
WZTi2T220kN1gMjdSbuPxT+IdkhP05pqDwxIyhSGDN2+TaB+xXdx7y/c2DKkPjWh
+FGMax4X+q2h1I5xs/fN6tkObU7qYe4R/dDgbafetFQPkBui1S7WHVeLbhJxVHKa
RAgWEKg2u1c0VgpaEGHqBtQEdm2b7PAIL7DIwbS++Z7gwGhM8Kj9KHkOA39LNC0u
+/jACrIqJ98ZyPkWwEtvXNzDBhEPZOuKCg/caN4Trv26Pzs/vFxmnisrN6Dqn00B
bbQzvDOfhSC8yEfjQpdA+G1bscsa+IaUCDbb7eNS4YVu8+UDm9k0u5byO2lfjgIT
VORd0b/VY1z9ht0dOrNFWaWam3VJovDJ7DoZn7CnZaz2XgbB6EhxGRIvbC0XhmVT
srqZ/PS8AD98dWQF5h3nMHsldmZ7picfJRiNrnlcpHCHAbcBfQbOadlkw3EpEaAf
Ah/bOBl+/V9vHtTvoapZFPtTNAJKv3+TW2MzrZ1GHmuROEh/tKiQkOEb8ZXFMomz
SwXzikEyZKpKjG1ZCAhARAUpD/dnRgtfwTP0FwiK/shJz3sXiB3QpyPr228zM2c1
8UwzbHTGYJ5cLj0L29+YspA68pzjdMsY7IZ5QJVv1jiH/FwP4JX/1jSy4OQr0iRv
InszgVyJ6KPlA4PRbTFWkHZyBC1sMWBxebwpAJvfXEjghBvkW6aXDe5NLVtcTcjk
43rbxYoC9OKs8D4lBbtvAr4z5gfGJlNjcSi6N9fTmNcH5Rg5lcG+LpMRsFNUIkBc
6fSiC2ukuyCI/6F2VX8olmDSPgOyYfbDxIaGQimQKpeIWnmpBvW3MhzgpN9QLB6X
S1LCHdq3amXAhMyldeOwvb7yk5OOwRHDPz+x/XrnZPqA4vNERAAvY87y3NJXyFOy
4Vm7Jc/3e3FhLuStVZcnx2ksv9gMG38Vq/mMBWDrFnyP7/5k11sHz6wTORO4ugWW
H6nbbOxXYT9Ac8dl5hVz8YoudimajucXyoWsczrDCoJbj21RZzAeib+2CbCdK4g+
I6PF9Lq4DXbd+McWusHrlUEGv10D/hxnMMeHRMcn5y8GgfbRPDblhdnFC0AjAwE5
8xnrVkoB3PtbnjyrnGFJyGoHb/tf3NJA1XhfK4kqDZI1cFWRq3llu0ZxC466s30K
uwQPcQ0udi2iaoKootxDw7QViQg+bZ7BtXgozaebQEMqTpmkK5QDFQmjB6qjP9o7
yG8OELC5rnAu7dNR+E2yr8GrxNTSIrwAQJu8RweVjsKpMccUImenBMEhh+a5ktkB
tP5zO8TnSCZ0oawdKQ5x3gClCkmYcGIEMhcYyTMwyuWMZcBCESQREFWOfQH1LzcE
8A6RY3sx9dpJNIqB08CpIR/tyO2X1zdTusT6dYk6i2Kxt7ekVigJU1lNivn3pEJ7
gTBgxVTPm6uqGpLZVnPIKlVluxKA3fLLid8+5F0BxG1dPRcAa5x1KeLMJLUc+8/O
Q4nc0FqBCZHs+Nd9Rc+O5Wm4OBd2UB0Y6/HzobAP2WveobY1z/UACnug4PmHIDWv
TS12gn03oY1B4pnBYtOAS30dCm2Pd6mcE43xvS7ae74wjavXu7tGSsNGfQWazeL3
s3uG6vz7MtuuB6YPVP75R3xOyhkaM4SrOVFk+Nlcuz3PZOITBQaIlJdmnMdki18N
fEf7rtnulF0Iv4qiUOVS25NqQiW/y/VT1DDcqLUmycbqkn8Z7jFMdTQ4WbHnPNy/
t4OqwegBxzF1ngM0Mu8mQOaZ4P4oWetO+djOsM5SBiRCzzXZRe9bA7QWfl8IrnXx
8txWpoLfGg+DjoDS9oSyVDnGq1DY309w62jrlsncZUGecORjx91G+RmZXJUgxkco
MFgt2NJhodNIsW0fuxwekd+ZxQIc55JAZzLPLi3epei9CzTCkOFjEjPqwtvohj2O
RRNErUUm1ZTZs43TVFvp0biLvNZIVnmmxarX3dZOJeesSYOSzMsuL2nhJz9YS5zn
PzgRbjoi739tVNSSFN/Qe8xKfxWLZAmOag9EE6IqPbzDm3YnRUzNuSPk7e54fYZ+
D/HH3D8dMPrVbdxRLyN2eXvYPnNtHu7buqcws16qkAKqWvsDB0D72tsRUuBBudJn
ByD1LnVE9wQFPxPdnXcmO3lYS6MvNDUa/RBLJ5ompR3IZn9l5/IvwmwzYJPar4Sp
XYqjbt1xnbE3FzoW3N4qaPWL6jldJt6SzAwhqDMvk2m9v1NCFAkqZG5TVfhmbZHo
YWDC7X/L18tuRLncKI2mcMX7azGx8Z1eYxts9EpTVkk1B6V9m01n5nREK/Y4u/6d
PsU0eWITVgcjj7ymG0tKK/QW71+Jh0BPLyiFOpJ7/AqpAPJ3HQzkUguHlxe5Ykoa
MGFuYIc0Kv5By98O+1hIyeM0DJNOKvVaixiP8pL6lj6tK4FuBwhSbrAlFR2Onekb
nsTfZho67ITpJUCsthv0tIgmlwo4SfOFeNUyPdbnOp7N/5YC0ulG4D5dMzl/Gl5n
ZZTlD0Q4cRbP+vfnTBEWY6lJn6TsrIjKgRfwCiw7DXYtaASleoad5Ne7nXkH53qr
v3hJat9DH+/qkGyXyJ6l4LSRqk9R1g6ermsyLRthXlLlmStOfKbJXquoAXZ7AyME
NZkHiG19x3msSeVwJ+aa3IMQgdYJQr30O+Yo10OWs+7/e/tHx8+SPbjweNdlXsRg
Pd/KbdxfTtcxaRZc89zYwCsKxBFJ5MGfr1ixtP2MT+4a0tDBB6b/h21a48+9Uci1
Ij7CkE31iv24VUYC0OQDCg4s+Ye8GD5D3hR6Yv73Brj49ETVyhGLjvaYh2OqHuiJ
juHn3ZUxHrFES1eBBGYCShGrECKytdDxm3bIP5gCXtJrVgAEVjYxmleBBHTQuOAj
zxHcM47ZaXiseEw2gT4lDc9MZYJ8FLbXb8CrzWyDUG/wZl1idOcovuhE/8laqYxr
VBDtPnnjeE2lIGg+EHHxND9xjb43+Kndy4wZ21n/WDunq90lz59n6fnHxh1eg7k6
9QCRLl9as+CGx1Cw+rqtL+81bBQRpT8s5YXSVltRagZXoooVK8fJRD4L0XOLknn8
BUfYW8NweNEoht6pUPm1lnooz1qyGrn9t2dE8OMgtZXj3IuVjl808P2pK3rQGZ4L
Lza8uo8WO5NVac4g/wMmBDGeTW0lMEwIPTFhuDD3WTjoPEp6xFqAnblgJLYs21mI
mBb4z1UMQN75+zHhQSGnVC1wbIDnc/n5fPrOn30BpQwkufZ6el837unejYYvZZfr
ZPrppHBEW0MzevPYwtHJB9HNxQv6hqhtJ88SK1Bv41yf/IAvJaO7dlMpjiv2O8Pi
ndqsQFa5WjNturI8ZifoGnxSJJ/rR1kdn+mvDQ0OEDgbtfS8XAYWW3RwOUTMU8TT
aOTKpwctuiDg/QoDNSaNQpJN502uvdjoMElp7NbWKofQwLbsSJL8jTCam1JLywVG
izf4r6zq4/gFTg4JRkLjSjqGvO3Dt2qwt6bFzkurUUf7u8na77SIHBjSmJgoum3q
1q1ueUq7pGxRWzY144kQh0mQbCn4D5irbkFaSrSnQL5eaUmXtoETfVNYR2o95zzA
aORHKl5JFUAyKqogICF8NPW83lhM21fQyYO3Vnav868tBli8/6TFmDyzR3IzftMs
CFE5H8cJ1G0m9awcujxfU6WUj2tWbgYzRzTKM0nO/7wey/hMS19R4qP2acC1cWBH
c1E66i/2EFKcf5zLlNxGSrDy6QedIAhc8CfDEtXU9vRjkkYj3h7UOxSM431t7UCW
0Wgm6adgjgPEXQOLc7DJDSVWh6kiV0WpNh6Sd2LqgWBZmD6vtwNe1SV/XJphUoN7
QH9xGJku+vOr2caYYvMgiWujW3Dhvr6kLYGIsMP++HieVez47NB1wUs0Fh5E3A71
C1OOj5IXH1fkBDDKpEiYsR76CtQH7GGP5gxo8gZdlbF1lYkiFAMbJzfFLJbQaNec
9sZNqsy00ILRYNcnuYHc2tunlCYZ42WA/OB+MVKmYUG8aEcsZ3aTBYuB/zxLp5Hm
9iHIchMSbdgDO/XEefVCYzDWHwEDB8usXloU4FfNpmz3kTNeT6q0IyRv+okvreGE
ueToDStA2E1pY+sgfaqbtWClDfu7uD7/zEHQIrhIu3+ZQQnQxFzfdyrR2g3yMp0p
TORtpgFv2JnP1eq/z6ZVjwm2BmEgxa1yqF0/iS4ycUlMft4i8uBWM8NxYojB2ZOh
Z016s9Kt+pbWSRkkb07IJA7SQ37ErOeRxscR0dZnVXGsPfFFn8h+mwcHLCIMBOKp
agbHevyviMzyXDNDbRJsL0Kf762eKjleE3RhMjQqGYIF7uLW6skF5h6Sf4ltbq67
gnJgx4wvE2Kpbsh6wqnFAFTjQYvEyxPpjwlxHPTvN9U7u2nBQAbCfxnIOvD0Gw2E
HxRizKsmeIyZ40ayM+bBOJioObbfQBU6THXWHnHzReeaRtSNMnvGnyMXnUmytyRP
1EK83vkIrVrxZ57jvt6eJj04/ccuko47KcUBh9/+ml6v+ix5yw0DHl/aKlezdxe3
JyUtIef1vsdONfVwFa2ky0VEFkCdQwSst1teqI/781Cq+29hVvDZDyUKNwamqvga
nzCIlulLsYC5W+1iDN0ufFjZ4fYBYZZO/+pSxPQV6NQHCQMjayJ6rOAgCL6VTB5z
6Q/9eQnDNwF/NPLair3d/5m8W0Jw6ZKMkvo1KwPvdLcZKBrhvFn1xALaYr3tuVta
qyR8D26+HrRlAag5T2UrI8JTmCsskfdoimbVZUln7AGKBrwCb70ANfrEmBC6R9ku
JCpNR+Z86ua9JUw+V0mFN2EnnR0oJ9SlIfyIzyZ9Rk2REhwRXHx25uePVVubPdF2
+uwnBGKylvcQfaSqm4zWEz+aAjKTWr1Yikf8d5ViE9H4Wl6piXhNzI6qiMMDa5IW
JAkzT5u/j2emx5kN8R72zoS+ysGKkp+ZytD2EzTNe1eiGEhvYpWqENmrbtCv/uxB
tmNs5rk1dzNv3MjfccbpWsUYfLcNg8FKyqEmeR7pej1kYoI1TbGPP/suZv1n3EaT
9FzEF17lNwNYIa44OsKElw+bT7d/fhvzY5K7rQE8gPYx+vnnlMP3qI/Q3tM/mKUW
yVPCsVC3AtYGUq1hDNPpjl4GzOLXWFr7NnGbqpBpr6chbZkrgn0VsDye5HKvQ1wP
e9iyoY/+WbbC2rbOLwfogg/GXQviqDR/39BhR6RkATX9+DvGqBJ3O4gQp651hwhw
nIMOJteC+/V033Nxl+i0PzPoiYumxKO5w+tN0x4T2SWlSmVPzSzM0+HuY5z1wZu+
xQTffp1VcxLutPM8dHgg3mc9WRVjB+XhDS6rTLL2hZkEw0t389uTCv9QJJl4za8S
8a0u28plHFcW3VBILrQmyxUP+OWWJrZ+hutw3MRJDv8Zeb0QDz1oqRUKVO0IzIRa
vIeOXFA91R+4kcWj6YySTtvGMxBvafj6koCJNeesBUnQ5Fz76N55WoaiwjdHIpgu
yrlfZW7gbA3JCXdlT1OvSmjUgW4hG0hQrbOfrr3W14uNSguLFYfrtGqaGRe/5ftg
uBYSkkr3lSMKp8QYui5GxjGPwGRFkxHhSjxl3ron+qnF9MJY4hbihESYeOsIn/jh
W6fRlWZmrRx6nSyXvxxcS6T0dnG6+pa1C63gqZEmY99Q91KzaZF80T7DiD8xagn3
TpyagrmelA/qjFRTDAEogb4bJYRAt0535ozS6O3iSk9srObcN13Kc18o7ldZpryq
WR/afApJKUYQRxrlji2qwfS1jfgyvRY8ltUrJCS36+o2Ua0D9VPSiILBgYBtw3MP
iNWU1OzMuR74krmyOaaDChcDiqG5NmDwEu/fVOwSGf25D4R31cSckz5k/ZJ1wV55
154bvA6ul1G8txitVxO8oInNVCr76O0xMpHP6STgN5kAzTrDH4VCeeZ+pso84yl/
FEYsaGL/VOSEEPfngj0WyfdtHk9oaHsqDng6FKGzhzxKPKj0LB6a4yV6DtrBY/0N
gZju0mIcMiulI/Q84D+Y7eJR5pVeyrr/0dt+v6GRyIYPGpHxNggQ8dTdSqrngyYe
NYCap83tKnPIGBtBV3Y8oOyWxeMj8JKuWdSFk9R3pbh+Gu9+oxq7//rbtQ/d1KIi
VVZNwpxvJ3rTWIwttj41CP5D6map+kdHoOiH3ugwg+xwD1zbA9lZilvhdLD4+amm
uvdB26bqW3QJN7daJQ42i7qSwsz6HoUDAKQo1sv/j5iM1NVfX+CIhYPk2z3cy8yy
Ph7fyAwydZxTPZUAQHLUjGE8x5SbeTwGA7b7RxYSI7t9Etx7ha5Tx1+LjzwRa63g
9tegsRK8p/u9Njj+tsgj7EOQ/zTBCBSGUuzCiN7YASElq5fls91IM3uaxBi9COrw
967iW76axDHvOwWZMneD0gE5cHN8wXOeT7S1Rla8clLHw9Ut/EEma96uMLEL2gd5
65gY1AmAKgQMKFxtDqlI8FGW7JPhjSXSg/DstTZHWaQL/1mkZ9LUgc0CbZI26Ine
1srWffiELhSCOzQYyGzI1bS0s2GfrSgvl42Teo+bb6R0LRBzvrQB8nk3znXo24oC
2Xa7sQlJsNO/spa1V6Rn4nlFugA2p82YDZl8bTNO+QoVudndwCR1UM9PhpikdC7H
nEy+ENJItjhpHUKkK2kFh6e9q6PnVfgBaJr+6A992FszA5dmcqBA3Gad+qGcCNne
qBuA7DOwsfDduoOzx2RqLgLLJZTY9/H5wYnbOPPDNS3aJjZ+FZ8LRGAd4PEgOMr4
YIMHsya5vzYLeM2RYlqIvKZSF5PcxoA4dcOIkLIM76F7HfoPZleh/27ceuyjBqQn
ssTE8DV9ctyfjYbvp8hQVaQSR+mpGJKbYNel3dztVSqQWtyPeop8AY6KBUQRLAmt
Z0Rr39dOWEJi4je8OdQmlbCIxI5hAvRW9NOEkC3uLkq5hHkvW5dTCGQhtjCVQMpv
9L7OZKzeHN5sMZKkmSryiUWI0AN30gExu+oQ247Ee8io3hHxxNcUJ/q90WMWa34R
qBnKCsNK8sfqwUiBennMUZc6XyGNBsKNIT+/yWNe3MOm8JQ1Yd/kPd9SEgNFuXGB
gGxZnQJaKilNFXtwvGKuZds+p5FjZJagK68YUYRJCT0vsuHwexSEkBOhgxBGyQ9i
zG0uEmWqcRy1Fp1YWMBeb5P7h52PsihhjAqIupV8VUkQaySBFOpKIOmRsUAY1//U
zAaYnsLiyzwd6i3TZy+EORS4nrrSdrGQyd79WzTh5uutI9ILEhiXCDbO+0xw2+oy
EXKknfnaI1lm49kSmEnyAGZ3UjItToELRU+6bXzV4vOeEMkp0ZI9glj10RCslWbC
uMM0ea5vszyE/IFDEO8yNDTCvOUMnkJ4SxEYqytvF/Q23D+NSP0b1fF2eF8xXjUo
adkcwe36Zt7ygOddEjfem8Cy1OacSVKNRQpmaV2sg1XrWSbaE9fPIqlkoY4mpz4Z
azR/twi2eJcx3eFZjWzW/x8XPfQr0A2eW29H+EmU/ageJMnSxl723XHej/wHI86Y
+HEhxoSbRRWku3jEqjjkGoFxo77ZUhwPZhPfIpldMHg9Fj4uUvDUk53ywldo2pxy
ubETTI1NYLt4L3BQYSLgUzY6Txxo0zyje8wcnFa+rlq6oJlgAV/X9jnu7mp/vQl1
GH7NqGDLO7eJaVWoGDqSLsp3gvZz0oiqgi9XZj3TD+SNL5iKpjWCHLMf8bfDkUdd
bCChljX1HlUsCNdlJgy2/rYs/tIEwVam0igSjzH5M/qxLP0S2L2YZQ/lpRXtMaS9
33e2mrTJKo3u9rUStjGjS67aFleXOU/k5XrXJKfKlnFgIVTj8fdwBMh9SvZ/bjT/
MNCr6qL7DttS/U7kHQskIt7CMUrFIijlRMgxkNZhraKsxixvemPj5h0rrcQERnmw
THloWI5rZ7YusktQxkKAJgAfRQ6DkGKxHO9kyIZQRoAGM1rVexJTQnSishSmAeR4
HbrXI2uRHshxs20KxUi0oBo7/T2Ib4KZeNsF35PmzbDW8Vtj7tsfiTD5qoxYNFo4
w7Kaambrt7XiWGsqs8PPfWVGYODaJ9vPDNq9ehsNyx7xBctU9O5NyXLvDGIqyyky
ga0WWQUMvnXC45hRreLB75Q+pJlrBwP0KHBGoVA2HwijkFxtV3/ks1RGmhsb7saS
74F5qdnqwnpZtcaBmmbkyiSzkFO6FiEriRyBmAF8ZfrEQgaL2FzZ4gMCTFUGRYLu
bQxjr9q3wjRIer2WGV80BXQFKFqMhSFTCIlTHV1q0dbqGwAI0qHsp2GDauOiuNGy
8sHLWcexCnOV7w/kffPm2wTwupQ0XrhjYM0eGrjZV/+PviPc9V+iJc0z9VQjFjfU
etnocNHZmQTzYpvi1KKd3rFoXWsagLrb3ZdtdL9YVnUqRVKh/zu8y06LlzuP/MFE
c3JJcTDaipT88m2nw0ooHORFqKLsOQ2M+wz0yxp1kyLoyseYW9nLRvuc1V4SEEHR
XkCTYHfQ6MDsfehEec9JzLLa/PcI0l1uz6GDym8uUPOcXW9Eqfv2AIkpAmHjSmrk
2tHaU7WISO2DdfQI/wTSZEAR7ZHynYZu2zWtxZvXIzmwytvYjVIUqCW2E0fQ5YXq
//pragma protect end_data_block
//pragma protect digest_block
0lnWj7KLT82FZ7gQ0RWG6rWo6X8=
//pragma protect end_digest_block
//pragma protect end_protected
