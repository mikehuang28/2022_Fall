`include "Usertype_FD.sv"

program automatic PATTERN_FD(input clk, INF.PATTERN_FD inf);
import usertype::*;



endprogram